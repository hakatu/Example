code gi do